* simple Inverter -ketan
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.param asn = 0.42*2 *0.15
.param pdn = 2*(0.42 + 2*0.15 )
.param wp = 0.84 + 0.42
.param asp = wp*2*0.15
.param pdp = 2*(wp + 2*0.15)
*.param rise_time =0
*.param fall_time =0

*the voltage sources:
Vdd vdd gnd DC 1.8
V1 in gnd pulse(0 1.8 0p 20p 20p 1n 2n)


Xnot1 in vdd gnd out not1   ; Inverter of single drive strength
Xnot2 out vdd gnd out1 not1

.subckt not1 a vdd vss z        ; subcircuit for inverter of single drive strength
xm01 z a vdd vdd sky130_fd_pr__pfet_01v8 l=0.15 w={wp}  as={asp} ad={asp}   ps={pdp} pd={pdp}
xm02 z a vss vss sky130_fd_pr__nfet_01v8 l=0.15 w=0.42 as={asn} ad={asn} ps={pdn} pd={pdn}
.ends

* simulation command for Time analysis:
.tran 1ps 10ns 0 1p
.measure tran rise_time TRIG v(out) VAL=0.36 RISE=1 TARG v(out) VAL=1.44 RISE=1     ; measure rise and fall times
.measure tran fall_time TRIG v(out) VAL=1.44 FALL=1 TARG v(out) VAL=0.36 FALL=1
.measure tran error_time PARAM='abs(rise_time - fall_time)'                         ; measure error time between rise and fall times
.measure tran error_percent PARAM='error_time*100/rise_time'                        ; measure error percentage between rise and fall times
.measure tran P_delay_TpHL TRIG v(in) VAL= 0.9 RISE=1 TARG v(out) VAL=0.9 FALL=1    ; measure propagation delay from input to output for high to low
.measure tran P_delay_TpLH TRIG v(in) VAL= 0.9 FALL=1 TARG v(out) VAl=0.9 RISE=1    ; measure propagation delay from input to output for low to high
.measure tran P_delay_avg PARAM='(P_delay_TpHL + P_delay_TpLH)/2'                   ; measure average propagation delay

.control
run
plot v(out) v(in)
.endc